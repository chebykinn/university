`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:38:30 10/24/2016 
// Design Name: 
// Module Name:    reader 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module reader(
    input CLK,
    input CS,
    input SDO,
    output [7:0] data
    );
	 
	 reg[7:0] data;


endmodule
